module vga_if (
  input clkIn,
  input rstIn,
  output [3:0] vgaROut,
  output [3:0] vgaGOut,
  output [3:0] vgaBOut,
  output vgaHsOut,
  output vgaVsOut
);

  wire rstW = ~rstIn;

  always @ (posedge rstW, posedge clkIn) begin
    if (rstW == 1) begin
    end

    else if (clkIn == 1) begin
    end
  end

endmodule

/* 
Design Notes

1. At each pixel clock (the main clock generated by the PLL), the horizontal counter increments.
Once the counter reaches the maximum horizontal count, there is going to be a blanking time, which
inclues a front porch section, followed by a sync pulse, followed by a back porch section. During 
the sync pulse section, the H-Sync signal will be low. Every other time, H-Sync will be high.

2. Once the horizontal counter reaches the maximum horizontal count, the vertical counter will
increment. Once the vertical counter reaches the maximum vertical count, there is going to be
a blanking time, which includes the same sections mentioned above. During the sync pulse
section, the V-Sync signal will be low. Every other time, V-Sync will be high.

3. During the duration on the blanking period, make sure that all outputs are 0.

4. 
*/
